module kbd_ipod_controller (
                            clk,
                            kbd_received_ascii_code,
                            reset_address,
                            play_pause,
                        
)